module InstructionMemory (
    input clk,
    input rst,
    input [31: 0] PC,
    output [31: 0] Instruction
);

reg [31:0] InstructionMemoryData [511: 0];

assign Instruction = InstructionMemoryData[PC[10:2]];

always @(posedge rst) begin
InstructionMemoryData[9'h0] <= 32'h00000000;
InstructionMemoryData[9'h1] <= 32'h00000000;
InstructionMemoryData[9'h2] <= 32'h00000000;
InstructionMemoryData[9'h3] <= 32'h20080004;
InstructionMemoryData[9'h4] <= 32'hac080000;
InstructionMemoryData[9'h5] <= 32'h20080000;
InstructionMemoryData[9'h6] <= 32'hac080004;
InstructionMemoryData[9'h7] <= 32'h20080008;
InstructionMemoryData[9'h8] <= 32'hac080008;
InstructionMemoryData[9'h9] <= 32'h2008ffff;
InstructionMemoryData[9'ha] <= 32'hac08000c;
InstructionMemoryData[9'hb] <= 32'h2008ffff;
InstructionMemoryData[9'hc] <= 32'hac080010;
InstructionMemoryData[9'hd] <= 32'h20080005;
InstructionMemoryData[9'he] <= 32'hac080084;
InstructionMemoryData[9'hf] <= 32'h20080000;
InstructionMemoryData[9'h10] <= 32'hac080088;
InstructionMemoryData[9'h11] <= 32'h20080002;
InstructionMemoryData[9'h12] <= 32'hac08008c;
InstructionMemoryData[9'h13] <= 32'h20080004;
InstructionMemoryData[9'h14] <= 32'hac080090;
InstructionMemoryData[9'h15] <= 32'h2008ffff;
InstructionMemoryData[9'h16] <= 32'hac080104;
InstructionMemoryData[9'h17] <= 32'h20080002;
InstructionMemoryData[9'h18] <= 32'hac080108;
InstructionMemoryData[9'h19] <= 32'h20080000;
InstructionMemoryData[9'h1a] <= 32'hac08010c;
InstructionMemoryData[9'h1b] <= 32'h20080001;
InstructionMemoryData[9'h1c] <= 32'hac080110;
InstructionMemoryData[9'h1d] <= 32'h2008ffff;
InstructionMemoryData[9'h1e] <= 32'hac080184;
InstructionMemoryData[9'h1f] <= 32'h20080004;
InstructionMemoryData[9'h20] <= 32'hac080188;
InstructionMemoryData[9'h21] <= 32'h20080001;
InstructionMemoryData[9'h22] <= 32'hac08018c;
InstructionMemoryData[9'h23] <= 32'h20080000;
InstructionMemoryData[9'h24] <= 32'hac080190;
InstructionMemoryData[9'h25] <= 32'h20080000;
InstructionMemoryData[9'h26] <= 32'h8d040000;
InstructionMemoryData[9'h27] <= 32'h21050004;
InstructionMemoryData[9'h28] <= 32'h20080640;
InstructionMemoryData[9'h29] <= 32'had000000;
InstructionMemoryData[9'h2a] <= 32'h21090004;
InstructionMemoryData[9'h2b] <= 32'h00042080;
InstructionMemoryData[9'h2c] <= 32'h00885020;
InstructionMemoryData[9'h2d] <= 32'h200bffff;
InstructionMemoryData[9'h2e] <= 32'h112a0003;
InstructionMemoryData[9'h2f] <= 32'had2b0000;
InstructionMemoryData[9'h30] <= 32'h21290004;
InstructionMemoryData[9'h31] <= 32'h0800002e;
InstructionMemoryData[9'h32] <= 32'h20110004;
InstructionMemoryData[9'h33] <= 32'h12240023;
InstructionMemoryData[9'h34] <= 32'h20120000;
InstructionMemoryData[9'h35] <= 32'h1244001f;
InstructionMemoryData[9'h36] <= 32'h20130000;
InstructionMemoryData[9'h37] <= 32'h1264001b;
InstructionMemoryData[9'h38] <= 32'h00126940;
InstructionMemoryData[9'h39] <= 32'h01b36820;
InstructionMemoryData[9'h3a] <= 32'h01127020;
InstructionMemoryData[9'h3b] <= 32'h8dcf0000;
InstructionMemoryData[9'h3c] <= 32'h00000000;
InstructionMemoryData[9'h3d] <= 32'h00000000;
InstructionMemoryData[9'h3e] <= 32'h2001ffff;
InstructionMemoryData[9'h3f] <= 32'h102f0011;
InstructionMemoryData[9'h40] <= 32'h00ad7020;
InstructionMemoryData[9'h41] <= 32'h8dd80000;
InstructionMemoryData[9'h42] <= 32'h00000000;
InstructionMemoryData[9'h43] <= 32'h00000000;
InstructionMemoryData[9'h44] <= 32'h2001ffff;
InstructionMemoryData[9'h45] <= 32'h1038000b;
InstructionMemoryData[9'h46] <= 32'h0113b020;
InstructionMemoryData[9'h47] <= 32'h8ed90000;
InstructionMemoryData[9'h48] <= 32'h00000000;
InstructionMemoryData[9'h49] <= 32'h00000000;
InstructionMemoryData[9'h4a] <= 32'h01f8a020;
InstructionMemoryData[9'h4b] <= 32'h2001ffff;
InstructionMemoryData[9'h4c] <= 32'h10390003;
InstructionMemoryData[9'h4d] <= 32'h0334a822;
InstructionMemoryData[9'h4e] <= 32'h1ea00001;
InstructionMemoryData[9'h4f] <= 32'h08000051;
InstructionMemoryData[9'h50] <= 32'haed40000;
InstructionMemoryData[9'h51] <= 32'h22730004;
InstructionMemoryData[9'h52] <= 32'h08000037;
InstructionMemoryData[9'h53] <= 32'h22520004;
InstructionMemoryData[9'h54] <= 32'h08000035;
InstructionMemoryData[9'h55] <= 32'h22310004;
InstructionMemoryData[9'h56] <= 32'h08000033;
InstructionMemoryData[9'h57] <= 32'h21090004;
InstructionMemoryData[9'h58] <= 32'h20020000;
InstructionMemoryData[9'h59] <= 32'h00885020;
InstructionMemoryData[9'h5a] <= 32'h112a0006;
InstructionMemoryData[9'h5b] <= 32'h8d2b0000;
InstructionMemoryData[9'h5c] <= 32'h00000000;
InstructionMemoryData[9'h5d] <= 32'h00000000;
InstructionMemoryData[9'h5e] <= 32'h004b1020;
InstructionMemoryData[9'h5f] <= 32'h21290004;
InstructionMemoryData[9'h60] <= 32'h0800005a;
InstructionMemoryData[9'h61] <= 32'h2408000f;
InstructionMemoryData[9'h62] <= 32'h2409000f;
InstructionMemoryData[9'h63] <= 32'h00094900;
InstructionMemoryData[9'h64] <= 32'h240a000f;
InstructionMemoryData[9'h65] <= 32'h000a5200;
InstructionMemoryData[9'h66] <= 32'h240b000f;
InstructionMemoryData[9'h67] <= 32'h000b5b00;
InstructionMemoryData[9'h68] <= 32'h00488024;
InstructionMemoryData[9'h69] <= 32'h00498824;
InstructionMemoryData[9'h6a] <= 32'h00118902;
InstructionMemoryData[9'h6b] <= 32'h004a9024;
InstructionMemoryData[9'h6c] <= 32'h00129202;
InstructionMemoryData[9'h6d] <= 32'h004b9824;
InstructionMemoryData[9'h6e] <= 32'h00139b02;
InstructionMemoryData[9'h6f] <= 32'h24080004;
InstructionMemoryData[9'h70] <= 32'h00084700;
InstructionMemoryData[9'h71] <= 32'h21080010;
InstructionMemoryData[9'h72] <= 32'h00102021;
InstructionMemoryData[9'h73] <= 32'h24050001;
InstructionMemoryData[9'h74] <= 32'h0c000083;
InstructionMemoryData[9'h75] <= 32'h0c0000e2;
InstructionMemoryData[9'h76] <= 32'h00112021;
InstructionMemoryData[9'h77] <= 32'h24050002;
InstructionMemoryData[9'h78] <= 32'h0c000083;
InstructionMemoryData[9'h79] <= 32'h0c0000e2;
InstructionMemoryData[9'h7a] <= 32'h00122021;
InstructionMemoryData[9'h7b] <= 32'h24050004;
InstructionMemoryData[9'h7c] <= 32'h0c000083;
InstructionMemoryData[9'h7d] <= 32'h0c0000e2;
InstructionMemoryData[9'h7e] <= 32'h00132021;
InstructionMemoryData[9'h7f] <= 32'h24050008;
InstructionMemoryData[9'h80] <= 32'h0c000083;
InstructionMemoryData[9'h81] <= 32'h0c0000e2;
InstructionMemoryData[9'h82] <= 32'h08000072;
InstructionMemoryData[9'h83] <= 32'h24190fe0;
InstructionMemoryData[9'h84] <= 32'h0325c820;
InstructionMemoryData[9'h85] <= 32'h20010001;
InstructionMemoryData[9'h86] <= 32'h10240009;
InstructionMemoryData[9'h87] <= 32'h20010004;
InstructionMemoryData[9'h88] <= 32'h10240007;
InstructionMemoryData[9'h89] <= 32'h2001000b;
InstructionMemoryData[9'h8a] <= 32'h10240005;
InstructionMemoryData[9'h8b] <= 32'h2001000c;
InstructionMemoryData[9'h8c] <= 32'h10240003;
InstructionMemoryData[9'h8d] <= 32'h2001000d;
InstructionMemoryData[9'h8e] <= 32'h10240001;
InstructionMemoryData[9'h8f] <= 32'h08000092;
InstructionMemoryData[9'h90] <= 32'h20010020;
InstructionMemoryData[9'h91] <= 32'h0321c822;
InstructionMemoryData[9'h92] <= 32'h20010005;
InstructionMemoryData[9'h93] <= 32'h1024000b;
InstructionMemoryData[9'h94] <= 32'h20010006;
InstructionMemoryData[9'h95] <= 32'h10240009;
InstructionMemoryData[9'h96] <= 32'h2001000b;
InstructionMemoryData[9'h97] <= 32'h10240007;
InstructionMemoryData[9'h98] <= 32'h2001000c;
InstructionMemoryData[9'h99] <= 32'h10240005;
InstructionMemoryData[9'h9a] <= 32'h2001000e;
InstructionMemoryData[9'h9b] <= 32'h10240003;
InstructionMemoryData[9'h9c] <= 32'h2001000f;
InstructionMemoryData[9'h9d] <= 32'h10240001;
InstructionMemoryData[9'h9e] <= 32'h080000a1;
InstructionMemoryData[9'h9f] <= 32'h20010040;
InstructionMemoryData[9'ha0] <= 32'h0321c822;
InstructionMemoryData[9'ha1] <= 32'h20010002;
InstructionMemoryData[9'ha2] <= 32'h10240007;
InstructionMemoryData[9'ha3] <= 32'h2001000c;
InstructionMemoryData[9'ha4] <= 32'h10240005;
InstructionMemoryData[9'ha5] <= 32'h2001000e;
InstructionMemoryData[9'ha6] <= 32'h10240003;
InstructionMemoryData[9'ha7] <= 32'h2001000f;
InstructionMemoryData[9'ha8] <= 32'h10240001;
InstructionMemoryData[9'ha9] <= 32'h080000ac;
InstructionMemoryData[9'haa] <= 32'h20010080;
InstructionMemoryData[9'hab] <= 32'h0321c822;
InstructionMemoryData[9'hac] <= 32'h20010001;
InstructionMemoryData[9'had] <= 32'h10240009;
InstructionMemoryData[9'hae] <= 32'h20010004;
InstructionMemoryData[9'haf] <= 32'h10240007;
InstructionMemoryData[9'hb0] <= 32'h20010007;
InstructionMemoryData[9'hb1] <= 32'h10240005;
InstructionMemoryData[9'hb2] <= 32'h2001000a;
InstructionMemoryData[9'hb3] <= 32'h10240003;
InstructionMemoryData[9'hb4] <= 32'h2001000f;
InstructionMemoryData[9'hb5] <= 32'h10240001;
InstructionMemoryData[9'hb6] <= 32'h080000b9;
InstructionMemoryData[9'hb7] <= 32'h20010100;
InstructionMemoryData[9'hb8] <= 32'h0321c822;
InstructionMemoryData[9'hb9] <= 32'h20010001;
InstructionMemoryData[9'hba] <= 32'h1024000b;
InstructionMemoryData[9'hbb] <= 32'h20010003;
InstructionMemoryData[9'hbc] <= 32'h10240009;
InstructionMemoryData[9'hbd] <= 32'h20010004;
InstructionMemoryData[9'hbe] <= 32'h10240007;
InstructionMemoryData[9'hbf] <= 32'h20010005;
InstructionMemoryData[9'hc0] <= 32'h10240005;
InstructionMemoryData[9'hc1] <= 32'h20010007;
InstructionMemoryData[9'hc2] <= 32'h10240003;
InstructionMemoryData[9'hc3] <= 32'h20010009;
InstructionMemoryData[9'hc4] <= 32'h10240001;
InstructionMemoryData[9'hc5] <= 32'h080000c8;
InstructionMemoryData[9'hc6] <= 32'h20010200;
InstructionMemoryData[9'hc7] <= 32'h0321c822;
InstructionMemoryData[9'hc8] <= 32'h20010001;
InstructionMemoryData[9'hc9] <= 32'h1024000b;
InstructionMemoryData[9'hca] <= 32'h20010002;
InstructionMemoryData[9'hcb] <= 32'h10240009;
InstructionMemoryData[9'hcc] <= 32'h20010003;
InstructionMemoryData[9'hcd] <= 32'h10240007;
InstructionMemoryData[9'hce] <= 32'h20010007;
InstructionMemoryData[9'hcf] <= 32'h10240005;
InstructionMemoryData[9'hd0] <= 32'h2001000c;
InstructionMemoryData[9'hd1] <= 32'h10240003;
InstructionMemoryData[9'hd2] <= 32'h2001000d;
InstructionMemoryData[9'hd3] <= 32'h10240001;
InstructionMemoryData[9'hd4] <= 32'h080000d7;
InstructionMemoryData[9'hd5] <= 32'h20010400;
InstructionMemoryData[9'hd6] <= 32'h0321c822;
InstructionMemoryData[9'hd7] <= 32'h20010000;
InstructionMemoryData[9'hd8] <= 32'h10240005;
InstructionMemoryData[9'hd9] <= 32'h20010001;
InstructionMemoryData[9'hda] <= 32'h10240003;
InstructionMemoryData[9'hdb] <= 32'h20010007;
InstructionMemoryData[9'hdc] <= 32'h10240001;
InstructionMemoryData[9'hdd] <= 32'h080000e0;
InstructionMemoryData[9'hde] <= 32'h20010800;
InstructionMemoryData[9'hdf] <= 32'h0321c822;
InstructionMemoryData[9'he0] <= 32'had190000;
InstructionMemoryData[9'he1] <= 32'h03e00008;
InstructionMemoryData[9'he2] <= 32'h2416b1e0;
InstructionMemoryData[9'he3] <= 32'h24174e20;
InstructionMemoryData[9'he4] <= 32'h12d70012;
InstructionMemoryData[9'he5] <= 32'h00000000;
InstructionMemoryData[9'he6] <= 32'h00000000;
InstructionMemoryData[9'he7] <= 32'h00000000;
InstructionMemoryData[9'he8] <= 32'h00000000;
InstructionMemoryData[9'he9] <= 32'h00000000;
InstructionMemoryData[9'hea] <= 32'h00000000;
InstructionMemoryData[9'heb] <= 32'h00000000;
InstructionMemoryData[9'hec] <= 32'h00000000;
InstructionMemoryData[9'hed] <= 32'h00000000;
InstructionMemoryData[9'hee] <= 32'h00000000;
InstructionMemoryData[9'hef] <= 32'h00000000;
InstructionMemoryData[9'hf0] <= 32'h00000000;
InstructionMemoryData[9'hf1] <= 32'h00000000;
InstructionMemoryData[9'hf2] <= 32'h00000000;
InstructionMemoryData[9'hf3] <= 32'h00000000;
InstructionMemoryData[9'hf4] <= 32'h00000000;
InstructionMemoryData[9'hf5] <= 32'h22d60001;
InstructionMemoryData[9'hf6] <= 32'h080000e4;
InstructionMemoryData[9'hf7] <= 32'h03e00008;
end


endmodule